//**********************************************************
// RV32I instructions
`define RV32I_NOP		32'b00000000000000000000000000010011
`define RV32I_LUI		32'b?????????????????????????0110111
`define RV32I_AUIPC		32'b?????????????????????????0010111
`define RV32I_JAL		32'b?????????????????????????1101111
`define RV32I_JALR		32'b?????????????????000?????1100111
`define RV32I_BEQ		32'b?????????????????000?????1100011
`define RV32I_BNE		32'b?????????????????001?????1100011
`define RV32I_BLT		32'b?????????????????100?????1100011
`define RV32I_BGE		32'b?????????????????101?????1100011
`define RV32I_BLTU		32'b?????????????????110?????1100011
`define RV32I_BGEU		32'b?????????????????111?????1100011
`define RV32I_LB		32'b?????????????????000?????0000011
`define RV32I_LH		32'b?????????????????001?????0000011
`define RV32I_LW		32'b?????????????????010?????0000011
`define RV32I_LBU		32'b?????????????????100?????0000011
`define RV32I_LHU		32'b?????????????????101?????0000011
`define RV32I_SB		32'b?????????????????000?????0100011
`define RV32I_SH		32'b?????????????????001?????0100011
`define RV32I_SW		32'b?????????????????010?????0100011
`define RV32I_ADDI		32'b?????????????????000?????0010011
`define RV32I_SLTI		32'b?????????????????010?????0010011
`define RV32I_SLTIU		32'b?????????????????011?????0010011
`define RV32I_XORI		32'b?????????????????100?????0010011
`define RV32I_ORI		32'b?????????????????110?????0010011
`define RV32I_ANDI		32'b?????????????????111?????0010011
`define RV32I_SLLI		32'b0000000??????????001?????0010011
`define RV32I_SRLI		32'b0000000??????????101?????0010011
`define RV32I_SRAI		32'b0100000??????????101?????0010011
`define RV32I_ADD		32'b0000000??????????000?????0110011
`define RV32I_SUB		32'b0100000??????????000?????0110011
`define RV32I_SLL		32'b0000000??????????001?????0110011
`define RV32I_SLT		32'b0000000??????????010?????0110011
`define RV32I_SLTU		32'b0000000??????????011?????0110011
`define RV32I_XOR		32'b0000000??????????100?????0110011
`define RV32I_SRL		32'b0000000??????????101?????0110011
`define RV32I_SRA		32'b0100000??????????101?????0110011
`define RV32I_OR		32'b0000000??????????110?????0110011
`define RV32I_AND		32'b0000000??????????111?????0110011
`define RV32I_FENCE		32'b?????????????????000?????0001111
`define RV32I_ECALL		32'b00000000000000000000000001110011
`define RV32I_EBREAK	32'b00000000000100000000000001110011

//**********************************************************
// RV32M instructions
`define RV32M_MUL		32'b0000001??????????000?????0110011
`define RV32M_MULH		32'b0000001??????????001?????0110011
`define RV32M_MULHSU	32'b0000001??????????010?????0110011
`define RV32M_MULHU		32'b0000001??????????011?????0110011
`define RV32M_DIV		32'b0000001??????????100?????0110011
`define RV32M_DIVU		32'b0000001??????????101?????0110011
`define RV32M_REM		32'b0000001??????????110?????0110011
`define RV32M_REMU		32'b0000001??????????111?????0110011

//**********************************************************
// RV32F instructions
`define RV32F_FLW		32'b?????????????????010?????0000111
`define RV32F_FSW		32'b?????????????????010?????0100111
`define RV32F_FMADD		32'b?????00??????????????????1000011
`define RV32F_FMSUB		32'b?????00??????????????????1000111
`define RV32F_FNMSUB	32'b?????00??????????????????1001011
`define RV32F_FNMADD	32'b?????00??????????????????1001111
`define RV32F_FADD		32'b0000000??????????????????1010011
`define RV32F_FSUB		32'b0000100??????????????????1010011
`define RV32F_FMUL		32'b0001000??????????????????1010011
`define RV32F_FDIV		32'b0001100??????????????????1010011
`define RV32F_FSQRT		32'b010110000000?????????????1010011
`define RV32F_FSGNJ		32'b0010000??????????000?????1010011
`define RV32F_FSGNJN	32'b0010000??????????001?????1010011
`define RV32F_FSGNJX	32'b0010000??????????010?????1010011
`define RV32F_FMIN		32'b0010100??????????000?????1010011
`define RV32F_FMAX		32'b0010100??????????001?????1010011
`define RV32F_FCVT_W_S	32'b110000000000?????????????1010011
`define RV32F_FCVT_WU_S	32'b110000000001?????????????1010011
`define RV32F_FMV_X_W	32'b111000000000?????000?????1010011
`define RV32F_FEQ_S		32'b1010000??????????010?????1010011
`define RV32F_FLT_S		32'b1010000??????????001?????1010011
`define RV32F_FLE_S		32'b1010000??????????000?????1010011
`define RV32F_FCLASS_S	32'b111000000000?????001?????1010011
`define RV32F_FCVT_S_W	32'b110100000000?????????????1010011
`define RV32F_FCVT_S_WU	32'b110100000001?????????????1010011
`define RV32F_FMV_W_X	32'b111100000000?????000?????1010011

//**********************************************************
// write back source
`define SEL_ALU			3'd0
`define SEL_MEM			3'd1
`define SEL_MUL			3'd2
`define SEL_DIV			3'd3
`define SEL_FPU			3'd4

//**********************************************************
// ALU operations
`define ALU_ADD			4'd0
`define ALU_SUB			4'd1
`define ALU_AND			4'd2
`define ALU_OR			4'd3
`define ALU_XOR			4'd4
`define ALU_SLL			4'd5
`define ALU_SRL			4'd6
`define ALU_SRA			4'd7
`define ALU_SEQ			4'd8
`define ALU_SNE			4'd9
`define ALU_SLT			4'd10
`define ALU_SLTU		4'd11
`define ALU_SGE			4'd12
`define ALU_SGEU		4'd13
`define ALU_INC			4'd14

//**********************************************************
// MEM operations
`define MEM_LB			3'd0
`define MEM_LBU			3'd1
`define MEM_LH			3'd2
`define MEM_LHU			3'd3
`define MEM_LW			3'd4
`define MEM_SB			3'd5
`define MEM_SH			3'd6
`define MEM_SW			3'd7

//**********************************************************
// MUL operations
`define UMULL			2'd0
`define UMULH			2'd1
`define SMULH			2'd2
`define SUMULH			2'd3

//**********************************************************
// DIV operations
`define UDIV			2'd0
`define SDIV			2'd1
`define UREM			2'd2
`define SREM			2'd3

//**********************************************************
// CSR operations
`define CSR_RW			2'd0
`define CSR_RS			2'd1
`define CSR_RC			2'd2

//**********************************************************
// CSR addresses
`define CSR_ADDR_MISA	12'h301

//**********************************************************
// reset vector
`define RESET_VEC		32'h00000000



